vsfg
